library verilog;
use verilog.vl_types.all;
entity orientacion_vlg_check_tst is
    port(
        clearcountdoblar: in     vl_logic;
        o0              : in     vl_logic;
        o1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end orientacion_vlg_check_tst;

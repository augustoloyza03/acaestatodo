library verilog;
use verilog.vl_types.all;
entity control3_vlg_vec_tst is
end control3_vlg_vec_tst;

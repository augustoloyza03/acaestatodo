library verilog;
use verilog.vl_types.all;
entity sensorlinea_vlg_check_tst is
    port(
        sensorlimpio    : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end sensorlinea_vlg_check_tst;

-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Dec 01 18:58:19 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY sensorlinea IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        sensorlinea : IN STD_LOGIC := '0';
        sensorlimpio : OUT STD_LOGIC
    );
END sensorlinea;

ARCHITECTURE BEHAVIOR OF sensorlinea IS
    TYPE type_fstate IS (blanco,blanco1,blanco2,blanco3,blanco4,blanco5,negro,negro1,negro2,negro3,negro4,negro5);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='0') THEN
            fstate <= blanco;
        ELSIF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,sensorlinea)
    BEGIN
        sensorlimpio <= '0';
        CASE fstate IS
            WHEN blanco =>
                IF ((sensorlinea = '1')) THEN
                    reg_fstate <= blanco;
                ELSIF ((sensorlinea = '0')) THEN
                    reg_fstate <= blanco1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= blanco;
                END IF;

                sensorlimpio <= '1';
            WHEN blanco1 =>
                reg_fstate <= blanco2;

                sensorlimpio <= '1';
            WHEN blanco2 =>
                reg_fstate <= blanco3;

                sensorlimpio <= '1';
            WHEN blanco3 =>
                reg_fstate <= blanco4;

                sensorlimpio <= '1';
            WHEN blanco4 =>
                reg_fstate <= blanco5;

                sensorlimpio <= '1';
            WHEN blanco5 =>
                IF ((sensorlinea = '0')) THEN
                    reg_fstate <= negro;
                ELSIF ((sensorlinea = '1')) THEN
                    reg_fstate <= blanco;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= blanco5;
                END IF;

                sensorlimpio <= '1';
            WHEN negro =>
                IF ((sensorlinea = '0')) THEN
                    reg_fstate <= negro;
                ELSIF ((sensorlinea = '1')) THEN
                    reg_fstate <= negro1;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= negro;
                END IF;

                sensorlimpio <= '0';
            WHEN negro1 =>
                reg_fstate <= negro2;

                sensorlimpio <= '0';
            WHEN negro2 =>
                reg_fstate <= negro3;

                sensorlimpio <= '0';
            WHEN negro3 =>
                reg_fstate <= negro4;

                sensorlimpio <= '0';
            WHEN negro4 =>
                reg_fstate <= negro5;

                sensorlimpio <= '0';
            WHEN negro5 =>
                IF ((sensorlinea = '1')) THEN
                    reg_fstate <= blanco;
                ELSIF ((sensorlinea = '0')) THEN
                    reg_fstate <= negro;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= negro5;
                END IF;

                sensorlimpio <= '0';
            WHEN OTHERS => 
                sensorlimpio <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
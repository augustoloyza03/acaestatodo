library verilog;
use verilog.vl_types.all;
entity nueva_orientacion_vlg_vec_tst is
end nueva_orientacion_vlg_vec_tst;

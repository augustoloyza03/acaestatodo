library verilog;
use verilog.vl_types.all;
entity avanzar_vlg_vec_tst is
end avanzar_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity sensorlinea_vlg_vec_tst is
end sensorlinea_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity orientacion_vlg_vec_tst is
end orientacion_vlg_vec_tst;

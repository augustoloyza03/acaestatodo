-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- Created on Mon Nov 11 15:15:26 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY avanzar IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SENSOR_D : IN STD_LOGIC_VECTOR(11 DOWNTO 0) := "000000000000";
        SENSOR_I : IN STD_LOGIC_VECTOR(11 DOWNTO 0) := "000000000000";
        SALIDA_I : OUT STD_LOGIC_VECTOR(2 DOWNTO 0); ---- primer bit velocidad los otros son de motor
        SALIDA_D : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		  led1, led2: out std_LOGIC
    );
END avanzar;

ARCHITECTURE BEHAVIOR OF avanzar IS
    TYPE type_state IS (ocioso,Avanzar,CORRECCION_D,CORRECION_I);
    SIGNAL state : type_state;
BEGIN

    PROCESS (state,reset,SENSOR_D,SENSOR_I)
    BEGIN
        IF (reset='0') THEN
            state <= ocioso;
          
       elsif (rising_edge(clock)) then
            CASE state IS
                WHEN Avanzar =>
                    IF ((SENSOR_D(11 DOWNTO 0) <= "001011101110") AND (SENSOR_I(11 DOWNTO 0) > "001011101110")) THEN
                        state <= CORRECCION_D;
								led1 <= '1';
								led2 <= '0';
                    ELSIF (((SENSOR_I(11 DOWNTO 0) <= "001011101110") AND (SENSOR_D(11 DOWNTO 0) > "001011101110"))) THEN
                        state <= CORRECION_I;
								led1 <= '0';
								led2 <= '1';
                    else
                        state <= Avanzar;
                    END IF;

                    SALIDA_I <= "110";

                    SALIDA_D <= "110";
                WHEN CORRECCION_D =>
                    IF (SENSOR_D(11 DOWNTO 0) >= "001011101110") THEN -- senSOR_D
                        state <= avanzar;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        state <= CORRECCION_D;
                    END IF;

                    SALIDA_D <= "110";

                    SALIDA_I <= "100";
                WHEN CORRECION_I => 
                    IF ( SENSOR_I(11 DOWNTO 0) >= "001011101110") THEN
                        state <= avanzar;
                   
                    ELSE
                        state <= CORRECION_I;
                    END IF;

                    SALIDA_D <= "100";

                    SALIDA_I <= "110";
              when ocioso =>
			       state <= avanzar;
					 SALIDA_I <= "100";
                SALIDA_D <= "100";
			
           END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;

library verilog;
use verilog.vl_types.all;
entity ubicacion_vlg_check_tst is
    port(
        clearcountdoblar: in     vl_logic;
        o0              : in     vl_logic;
        o1              : in     vl_logic;
        p0              : in     vl_logic;
        p1              : in     vl_logic;
        p2              : in     vl_logic;
        p3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ubicacion_vlg_check_tst;

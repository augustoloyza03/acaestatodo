library verilog;
use verilog.vl_types.all;
entity nueva_orientacion_vlg_check_tst is
    port(
        NO0             : in     vl_logic;
        NO1             : in     vl_logic;
        S0              : in     vl_logic;
        S1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end nueva_orientacion_vlg_check_tst;
